
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity tb_rowdecode is
    port (
        clk : in std_logic;
        rnd : in std_logic;
        rdy : out std_logic
    );
end entity tb_rowdecode;

architecture behavioral of tb_rowdecode is
signal rdy0 : std_logic;
signal row0 : std_logic_vector(13 downto 0);
signal rdy1 : std_logic;
signal row1 : std_logic_vector(13 downto 0);
signal rdy2 : std_logic;
signal row2 : std_logic_vector(13 downto 0);
signal rdy3 : std_logic;
signal row3 : std_logic_vector(13 downto 0);
signal rdy4 : std_logic;
signal row4 : std_logic_vector(13 downto 0);
signal rdy5 : std_logic;
signal row5 : std_logic_vector(13 downto 0);
signal rdy6 : std_logic;
signal row6 : std_logic_vector(13 downto 0);
signal rdy7 : std_logic;
signal row7 : std_logic_vector(13 downto 0);
signal rdy8 : std_logic;
signal row8 : std_logic_vector(13 downto 0);
signal rdy9 : std_logic;
signal row9 : std_logic_vector(13 downto 0);
signal rdy10 : std_logic;
signal row10 : std_logic_vector(13 downto 0);
signal rdy11 : std_logic;
signal row11 : std_logic_vector(13 downto 0);
signal rdy12 : std_logic;
signal row12 : std_logic_vector(13 downto 0);
signal rdy13 : std_logic;
signal row13 : std_logic_vector(13 downto 0);
signal rdy14 : std_logic;
signal row14 : std_logic_vector(13 downto 0);
signal rdy15 : std_logic;
signal row15 : std_logic_vector(13 downto 0);
signal rdy16 : std_logic;
signal row16 : std_logic_vector(13 downto 0);
signal rdy17 : std_logic;
signal row17 : std_logic_vector(13 downto 0);
signal rdy18 : std_logic;
signal row18 : std_logic_vector(13 downto 0);
signal rdy19 : std_logic;
signal row19 : std_logic_vector(13 downto 0);
signal rdy20 : std_logic;
signal row20 : std_logic_vector(13 downto 0);
signal rdy21 : std_logic;
signal row21 : std_logic_vector(13 downto 0);
signal rdy22 : std_logic;
signal row22 : std_logic_vector(13 downto 0);
signal rdy23 : std_logic;
signal row23 : std_logic_vector(13 downto 0);
signal rdy24 : std_logic;
signal row24 : std_logic_vector(13 downto 0);
signal rdy25 : std_logic;
signal row25 : std_logic_vector(13 downto 0);
signal rdy26 : std_logic;
signal row26 : std_logic_vector(13 downto 0);
signal rdy27 : std_logic;
signal row27 : std_logic_vector(13 downto 0);
signal rdy28 : std_logic;
signal row28 : std_logic_vector(13 downto 0);
signal rdy29 : std_logic;
signal row29 : std_logic_vector(13 downto 0);
signal rdy30 : std_logic;
signal row30 : std_logic_vector(13 downto 0);
signal rdy31 : std_logic;
signal row31 : std_logic_vector(13 downto 0);
signal rdy32 : std_logic;
signal row32 : std_logic_vector(13 downto 0);
signal rdy33 : std_logic;
signal row33 : std_logic_vector(13 downto 0);
signal rdy34 : std_logic;
signal row34 : std_logic_vector(13 downto 0);
signal rdy35 : std_logic;
signal row35 : std_logic_vector(13 downto 0);
signal rdy36 : std_logic;
signal row36 : std_logic_vector(13 downto 0);
signal rdy37 : std_logic;
signal row37 : std_logic_vector(13 downto 0);
signal rdy38 : std_logic;
signal row38 : std_logic_vector(13 downto 0);
signal rdy39 : std_logic;
signal row39 : std_logic_vector(13 downto 0);
signal rdy40 : std_logic;
signal row40 : std_logic_vector(13 downto 0);
signal rdy41 : std_logic;
signal row41 : std_logic_vector(13 downto 0);
signal rdy42 : std_logic;
signal row42 : std_logic_vector(13 downto 0);
signal rdy43 : std_logic;
signal row43 : std_logic_vector(13 downto 0);
signal rdy44 : std_logic;
signal row44 : std_logic_vector(13 downto 0);
signal rdy45 : std_logic;
signal row45 : std_logic_vector(13 downto 0);
signal rdy46 : std_logic;
signal row46 : std_logic_vector(13 downto 0);
signal rdy47 : std_logic;
signal row47 : std_logic_vector(13 downto 0);
signal rdy48 : std_logic;
signal row48 : std_logic_vector(13 downto 0);
signal rdy49 : std_logic;
signal row49 : std_logic_vector(13 downto 0);
signal rdy50 : std_logic;
signal row50 : std_logic_vector(13 downto 0);
signal rdy51 : std_logic;
signal row51 : std_logic_vector(13 downto 0);
signal rdy52 : std_logic;
signal row52 : std_logic_vector(13 downto 0);
signal rdy53 : std_logic;
signal row53 : std_logic_vector(13 downto 0);
signal rdy54 : std_logic;
signal row54 : std_logic_vector(13 downto 0);
signal rdy55 : std_logic;
signal row55 : std_logic_vector(13 downto 0);
signal rdy56 : std_logic;
signal row56 : std_logic_vector(13 downto 0);
signal rdy57 : std_logic;
signal row57 : std_logic_vector(13 downto 0);
signal rdy58 : std_logic;
signal row58 : std_logic_vector(13 downto 0);
signal rdy59 : std_logic;
signal row59 : std_logic_vector(13 downto 0);
signal rdy60 : std_logic;
signal row60 : std_logic_vector(13 downto 0);
signal rdy61 : std_logic;
signal row61 : std_logic_vector(13 downto 0);
signal rdy62 : std_logic;
signal row62 : std_logic_vector(13 downto 0);
signal rdy63 : std_logic;
signal row63 : std_logic_vector(13 downto 0);
signal rdy64 : std_logic;
signal row64 : std_logic_vector(13 downto 0);
signal rdy65 : std_logic;
signal row65 : std_logic_vector(13 downto 0);
signal rdy66 : std_logic;
signal row66 : std_logic_vector(13 downto 0);
signal rdy67 : std_logic;
signal row67 : std_logic_vector(13 downto 0);
signal rdy68 : std_logic;
signal row68 : std_logic_vector(13 downto 0);
signal rdy69 : std_logic;
signal row69 : std_logic_vector(13 downto 0);
signal rdy70 : std_logic;
signal row70 : std_logic_vector(13 downto 0);
signal rdy71 : std_logic;
signal row71 : std_logic_vector(13 downto 0);
signal rdy72 : std_logic;
signal row72 : std_logic_vector(13 downto 0);
signal rdy73 : std_logic;
signal row73 : std_logic_vector(13 downto 0);
signal rdy74 : std_logic;
signal row74 : std_logic_vector(13 downto 0);
signal rdy75 : std_logic;
signal row75 : std_logic_vector(13 downto 0);
signal rdy76 : std_logic;
signal row76 : std_logic_vector(13 downto 0);
signal rdy77 : std_logic;
signal row77 : std_logic_vector(13 downto 0);
signal rdy78 : std_logic;
signal row78 : std_logic_vector(13 downto 0);
signal rdy79 : std_logic;
signal row79 : std_logic_vector(13 downto 0);
signal rdy80 : std_logic;
signal row80 : std_logic_vector(13 downto 0);
signal rdy81 : std_logic;
signal row81 : std_logic_vector(13 downto 0);
signal rdy82 : std_logic;
signal row82 : std_logic_vector(13 downto 0);
signal rdy83 : std_logic;
signal row83 : std_logic_vector(13 downto 0);
signal rdy84 : std_logic;
signal row84 : std_logic_vector(13 downto 0);
signal rdy85 : std_logic;
signal row85 : std_logic_vector(13 downto 0);
signal rdy86 : std_logic;
signal row86 : std_logic_vector(13 downto 0);
signal rdy87 : std_logic;
signal row87 : std_logic_vector(13 downto 0);
signal rdy88 : std_logic;
signal row88 : std_logic_vector(13 downto 0);
signal rdy89 : std_logic;
signal row89 : std_logic_vector(13 downto 0);
signal rdy90 : std_logic;
signal row90 : std_logic_vector(13 downto 0);
signal rdy91 : std_logic;
signal row91 : std_logic_vector(13 downto 0);
signal rdy92 : std_logic;
signal row92 : std_logic_vector(13 downto 0);
signal rdy93 : std_logic;
signal row93 : std_logic_vector(13 downto 0);
signal rdy94 : std_logic;
signal row94 : std_logic_vector(13 downto 0);
signal rdy95 : std_logic;
signal row95 : std_logic_vector(13 downto 0);
signal rdy96 : std_logic;
signal row96 : std_logic_vector(13 downto 0);
signal rdy97 : std_logic;
signal row97 : std_logic_vector(13 downto 0);
signal rdy98 : std_logic;
signal row98 : std_logic_vector(13 downto 0);
signal rdy99 : std_logic;
signal row99 : std_logic_vector(13 downto 0);
signal buf: std_logic_vector(114 downto 0);
signal clk_bufg: std_logic;

begin  -- architecture behavioral


--BUFG:GeneralClockBuffer
--UltraScale
--XilinxHDLLanguageTemplate,version2018.1
BUFG_inst : BUFG
port map(
        O=>clk_bufg,  --1-bitoutput:Clockoutput
        I=>clk        --1-bitinput:Clockinput
    );
--EndofBUFG_instinstantiation


rowdecoder0: entity work.rowdecode
    port map (
        row => row0,
        clk => clk_bufg,
        rdy => rdy0
        );


rowdecoder1: entity work.rowdecode
    port map (
        row => row1,
        clk => clk_bufg,
        rdy => rdy1
        );


rowdecoder2: entity work.rowdecode
    port map (
        row => row2,
        clk => clk_bufg,
        rdy => rdy2
        );


rowdecoder3: entity work.rowdecode
    port map (
        row => row3,
        clk => clk_bufg,
        rdy => rdy3
        );


rowdecoder4: entity work.rowdecode
    port map (
        row => row4,
        clk => clk_bufg,
        rdy => rdy4
        );


rowdecoder5: entity work.rowdecode
    port map (
        row => row5,
        clk => clk_bufg,
        rdy => rdy5
        );


rowdecoder6: entity work.rowdecode
    port map (
        row => row6,
        clk => clk_bufg,
        rdy => rdy6
        );


rowdecoder7: entity work.rowdecode
    port map (
        row => row7,
        clk => clk_bufg,
        rdy => rdy7
        );


rowdecoder8: entity work.rowdecode
    port map (
        row => row8,
        clk => clk_bufg,
        rdy => rdy8
        );


rowdecoder9: entity work.rowdecode
    port map (
        row => row9,
        clk => clk_bufg,
        rdy => rdy9
        );


rowdecoder10: entity work.rowdecode
    port map (
        row => row10,
        clk => clk_bufg,
        rdy => rdy10
        );


rowdecoder11: entity work.rowdecode
    port map (
        row => row11,
        clk => clk_bufg,
        rdy => rdy11
        );


rowdecoder12: entity work.rowdecode
    port map (
        row => row12,
        clk => clk_bufg,
        rdy => rdy12
        );


rowdecoder13: entity work.rowdecode
    port map (
        row => row13,
        clk => clk_bufg,
        rdy => rdy13
        );


rowdecoder14: entity work.rowdecode
    port map (
        row => row14,
        clk => clk_bufg,
        rdy => rdy14
        );


rowdecoder15: entity work.rowdecode
    port map (
        row => row15,
        clk => clk_bufg,
        rdy => rdy15
        );


rowdecoder16: entity work.rowdecode
    port map (
        row => row16,
        clk => clk_bufg,
        rdy => rdy16
        );


rowdecoder17: entity work.rowdecode
    port map (
        row => row17,
        clk => clk_bufg,
        rdy => rdy17
        );


rowdecoder18: entity work.rowdecode
    port map (
        row => row18,
        clk => clk_bufg,
        rdy => rdy18
        );


rowdecoder19: entity work.rowdecode
    port map (
        row => row19,
        clk => clk_bufg,
        rdy => rdy19
        );


rowdecoder20: entity work.rowdecode
    port map (
        row => row20,
        clk => clk_bufg,
        rdy => rdy20
        );


rowdecoder21: entity work.rowdecode
    port map (
        row => row21,
        clk => clk_bufg,
        rdy => rdy21
        );


rowdecoder22: entity work.rowdecode
    port map (
        row => row22,
        clk => clk_bufg,
        rdy => rdy22
        );


rowdecoder23: entity work.rowdecode
    port map (
        row => row23,
        clk => clk_bufg,
        rdy => rdy23
        );


rowdecoder24: entity work.rowdecode
    port map (
        row => row24,
        clk => clk_bufg,
        rdy => rdy24
        );


rowdecoder25: entity work.rowdecode
    port map (
        row => row25,
        clk => clk_bufg,
        rdy => rdy25
        );


rowdecoder26: entity work.rowdecode
    port map (
        row => row26,
        clk => clk_bufg,
        rdy => rdy26
        );


rowdecoder27: entity work.rowdecode
    port map (
        row => row27,
        clk => clk_bufg,
        rdy => rdy27
        );


rowdecoder28: entity work.rowdecode
    port map (
        row => row28,
        clk => clk_bufg,
        rdy => rdy28
        );


rowdecoder29: entity work.rowdecode
    port map (
        row => row29,
        clk => clk_bufg,
        rdy => rdy29
        );


rowdecoder30: entity work.rowdecode
    port map (
        row => row30,
        clk => clk_bufg,
        rdy => rdy30
        );


rowdecoder31: entity work.rowdecode
    port map (
        row => row31,
        clk => clk_bufg,
        rdy => rdy31
        );


rowdecoder32: entity work.rowdecode
    port map (
        row => row32,
        clk => clk_bufg,
        rdy => rdy32
        );


rowdecoder33: entity work.rowdecode
    port map (
        row => row33,
        clk => clk_bufg,
        rdy => rdy33
        );


rowdecoder34: entity work.rowdecode
    port map (
        row => row34,
        clk => clk_bufg,
        rdy => rdy34
        );


rowdecoder35: entity work.rowdecode
    port map (
        row => row35,
        clk => clk_bufg,
        rdy => rdy35
        );


rowdecoder36: entity work.rowdecode
    port map (
        row => row36,
        clk => clk_bufg,
        rdy => rdy36
        );


rowdecoder37: entity work.rowdecode
    port map (
        row => row37,
        clk => clk_bufg,
        rdy => rdy37
        );


rowdecoder38: entity work.rowdecode
    port map (
        row => row38,
        clk => clk_bufg,
        rdy => rdy38
        );


rowdecoder39: entity work.rowdecode
    port map (
        row => row39,
        clk => clk_bufg,
        rdy => rdy39
        );


rowdecoder40: entity work.rowdecode
    port map (
        row => row40,
        clk => clk_bufg,
        rdy => rdy40
        );


rowdecoder41: entity work.rowdecode
    port map (
        row => row41,
        clk => clk_bufg,
        rdy => rdy41
        );


rowdecoder42: entity work.rowdecode
    port map (
        row => row42,
        clk => clk_bufg,
        rdy => rdy42
        );


rowdecoder43: entity work.rowdecode
    port map (
        row => row43,
        clk => clk_bufg,
        rdy => rdy43
        );


rowdecoder44: entity work.rowdecode
    port map (
        row => row44,
        clk => clk_bufg,
        rdy => rdy44
        );


rowdecoder45: entity work.rowdecode
    port map (
        row => row45,
        clk => clk_bufg,
        rdy => rdy45
        );


rowdecoder46: entity work.rowdecode
    port map (
        row => row46,
        clk => clk_bufg,
        rdy => rdy46
        );


rowdecoder47: entity work.rowdecode
    port map (
        row => row47,
        clk => clk_bufg,
        rdy => rdy47
        );


rowdecoder48: entity work.rowdecode
    port map (
        row => row48,
        clk => clk_bufg,
        rdy => rdy48
        );


rowdecoder49: entity work.rowdecode
    port map (
        row => row49,
        clk => clk_bufg,
        rdy => rdy49
        );


rowdecoder50: entity work.rowdecode
    port map (
        row => row50,
        clk => clk_bufg,
        rdy => rdy50
        );


rowdecoder51: entity work.rowdecode
    port map (
        row => row51,
        clk => clk_bufg,
        rdy => rdy51
        );


rowdecoder52: entity work.rowdecode
    port map (
        row => row52,
        clk => clk_bufg,
        rdy => rdy52
        );


rowdecoder53: entity work.rowdecode
    port map (
        row => row53,
        clk => clk_bufg,
        rdy => rdy53
        );


rowdecoder54: entity work.rowdecode
    port map (
        row => row54,
        clk => clk_bufg,
        rdy => rdy54
        );


rowdecoder55: entity work.rowdecode
    port map (
        row => row55,
        clk => clk_bufg,
        rdy => rdy55
        );


rowdecoder56: entity work.rowdecode
    port map (
        row => row56,
        clk => clk_bufg,
        rdy => rdy56
        );


rowdecoder57: entity work.rowdecode
    port map (
        row => row57,
        clk => clk_bufg,
        rdy => rdy57
        );


rowdecoder58: entity work.rowdecode
    port map (
        row => row58,
        clk => clk_bufg,
        rdy => rdy58
        );


rowdecoder59: entity work.rowdecode
    port map (
        row => row59,
        clk => clk_bufg,
        rdy => rdy59
        );


rowdecoder60: entity work.rowdecode
    port map (
        row => row60,
        clk => clk_bufg,
        rdy => rdy60
        );


rowdecoder61: entity work.rowdecode
    port map (
        row => row61,
        clk => clk_bufg,
        rdy => rdy61
        );


rowdecoder62: entity work.rowdecode
    port map (
        row => row62,
        clk => clk_bufg,
        rdy => rdy62
        );


rowdecoder63: entity work.rowdecode
    port map (
        row => row63,
        clk => clk_bufg,
        rdy => rdy63
        );


rowdecoder64: entity work.rowdecode
    port map (
        row => row64,
        clk => clk_bufg,
        rdy => rdy64
        );


rowdecoder65: entity work.rowdecode
    port map (
        row => row65,
        clk => clk_bufg,
        rdy => rdy65
        );


rowdecoder66: entity work.rowdecode
    port map (
        row => row66,
        clk => clk_bufg,
        rdy => rdy66
        );


rowdecoder67: entity work.rowdecode
    port map (
        row => row67,
        clk => clk_bufg,
        rdy => rdy67
        );


rowdecoder68: entity work.rowdecode
    port map (
        row => row68,
        clk => clk_bufg,
        rdy => rdy68
        );


rowdecoder69: entity work.rowdecode
    port map (
        row => row69,
        clk => clk_bufg,
        rdy => rdy69
        );


rowdecoder70: entity work.rowdecode
    port map (
        row => row70,
        clk => clk_bufg,
        rdy => rdy70
        );


rowdecoder71: entity work.rowdecode
    port map (
        row => row71,
        clk => clk_bufg,
        rdy => rdy71
        );


rowdecoder72: entity work.rowdecode
    port map (
        row => row72,
        clk => clk_bufg,
        rdy => rdy72
        );


rowdecoder73: entity work.rowdecode
    port map (
        row => row73,
        clk => clk_bufg,
        rdy => rdy73
        );


rowdecoder74: entity work.rowdecode
    port map (
        row => row74,
        clk => clk_bufg,
        rdy => rdy74
        );


rowdecoder75: entity work.rowdecode
    port map (
        row => row75,
        clk => clk_bufg,
        rdy => rdy75
        );


rowdecoder76: entity work.rowdecode
    port map (
        row => row76,
        clk => clk_bufg,
        rdy => rdy76
        );


rowdecoder77: entity work.rowdecode
    port map (
        row => row77,
        clk => clk_bufg,
        rdy => rdy77
        );


rowdecoder78: entity work.rowdecode
    port map (
        row => row78,
        clk => clk_bufg,
        rdy => rdy78
        );


rowdecoder79: entity work.rowdecode
    port map (
        row => row79,
        clk => clk_bufg,
        rdy => rdy79
        );


rowdecoder80: entity work.rowdecode
    port map (
        row => row80,
        clk => clk_bufg,
        rdy => rdy80
        );


rowdecoder81: entity work.rowdecode
    port map (
        row => row81,
        clk => clk_bufg,
        rdy => rdy81
        );


rowdecoder82: entity work.rowdecode
    port map (
        row => row82,
        clk => clk_bufg,
        rdy => rdy82
        );


rowdecoder83: entity work.rowdecode
    port map (
        row => row83,
        clk => clk_bufg,
        rdy => rdy83
        );


rowdecoder84: entity work.rowdecode
    port map (
        row => row84,
        clk => clk_bufg,
        rdy => rdy84
        );


rowdecoder85: entity work.rowdecode
    port map (
        row => row85,
        clk => clk_bufg,
        rdy => rdy85
        );


rowdecoder86: entity work.rowdecode
    port map (
        row => row86,
        clk => clk_bufg,
        rdy => rdy86
        );


rowdecoder87: entity work.rowdecode
    port map (
        row => row87,
        clk => clk_bufg,
        rdy => rdy87
        );


rowdecoder88: entity work.rowdecode
    port map (
        row => row88,
        clk => clk_bufg,
        rdy => rdy88
        );


rowdecoder89: entity work.rowdecode
    port map (
        row => row89,
        clk => clk_bufg,
        rdy => rdy89
        );


rowdecoder90: entity work.rowdecode
    port map (
        row => row90,
        clk => clk_bufg,
        rdy => rdy90
        );


rowdecoder91: entity work.rowdecode
    port map (
        row => row91,
        clk => clk_bufg,
        rdy => rdy91
        );


rowdecoder92: entity work.rowdecode
    port map (
        row => row92,
        clk => clk_bufg,
        rdy => rdy92
        );


rowdecoder93: entity work.rowdecode
    port map (
        row => row93,
        clk => clk_bufg,
        rdy => rdy93
        );


rowdecoder94: entity work.rowdecode
    port map (
        row => row94,
        clk => clk_bufg,
        rdy => rdy94
        );


rowdecoder95: entity work.rowdecode
    port map (
        row => row95,
        clk => clk_bufg,
        rdy => rdy95
        );


rowdecoder96: entity work.rowdecode
    port map (
        row => row96,
        clk => clk_bufg,
        rdy => rdy96
        );


rowdecoder97: entity work.rowdecode
    port map (
        row => row97,
        clk => clk_bufg,
        rdy => rdy97
        );


rowdecoder98: entity work.rowdecode
    port map (
        row => row98,
        clk => clk_bufg,
        rdy => rdy98
        );


rowdecoder99: entity work.rowdecode
    port map (
        row => row99,
        clk => clk_bufg,
        rdy => rdy99
        );


dummy_proc:process(clk, rnd) begin
    if rising_edge(clk) then
        rdy <= rdy0 xor rdy1 xor rdy2 xor rdy3 xor rdy4 xor rdy5 xor rdy6 xor rdy7 xor rdy8 xor rdy9 xor rdy10 xor rdy11 xor rdy12 xor rdy13 xor rdy14 xor rdy15 xor rdy16 xor rdy17 xor rdy18 xor rdy19 xor rdy20 xor rdy21 xor rdy22 xor rdy23 xor rdy24 xor rdy25 xor rdy26 xor rdy27 xor rdy28 xor rdy29 xor rdy30 xor rdy31 xor rdy32 xor rdy33 xor rdy34 xor rdy35 xor rdy36 xor rdy37 xor rdy38 xor rdy39 xor rdy40 xor rdy41 xor rdy42 xor rdy43 xor rdy44 xor rdy45 xor rdy46 xor rdy47 xor rdy48 xor rdy49 xor rdy50 xor rdy51 xor rdy52 xor rdy53 xor rdy54 xor rdy55 xor rdy56 xor rdy57 xor rdy58 xor rdy59 xor rdy60 xor rdy61 xor rdy62 xor rdy63 xor rdy64 xor rdy65 xor rdy66 xor rdy67 xor rdy68 xor rdy69 xor rdy70 xor rdy71 xor rdy72 xor rdy73 xor rdy74 xor rdy75 xor rdy76 xor rdy77 xor rdy78 xor rdy79 xor rdy80 xor rdy81 xor rdy82 xor rdy83 xor rdy84 xor rdy85 xor rdy86 xor rdy87 xor rdy88 xor rdy89 xor rdy90 xor rdy91 xor rdy92 xor rdy93 xor rdy94 xor rdy95 xor rdy96 xor rdy97 xor rdy98 xor rdy99 xor rnd;

buf <= std_logic_vector(shift_left(unsigned(buf), 1));
buf(29) <= rnd;

row0 <= buf(13 downto 0);
row1 <= buf(14 downto 1);
row2 <= buf(15 downto 2);
row3 <= buf(16 downto 3);
row4 <= buf(17 downto 4);
row5 <= buf(18 downto 5);
row6 <= buf(19 downto 6);
row7 <= buf(20 downto 7);
row8 <= buf(21 downto 8);
row9 <= buf(22 downto 9);
row10 <= buf(23 downto 10);
row11 <= buf(24 downto 11);
row12 <= buf(25 downto 12);
row13 <= buf(26 downto 13);
row14 <= buf(27 downto 14);
row15 <= buf(28 downto 15);
row16 <= buf(29 downto 16);
row17 <= buf(30 downto 17);
row18 <= buf(31 downto 18);
row19 <= buf(32 downto 19);
row20 <= buf(33 downto 20);
row21 <= buf(34 downto 21);
row22 <= buf(35 downto 22);
row23 <= buf(36 downto 23);
row24 <= buf(37 downto 24);
row25 <= buf(38 downto 25);
row26 <= buf(39 downto 26);
row27 <= buf(40 downto 27);
row28 <= buf(41 downto 28);
row29 <= buf(42 downto 29);
row30 <= buf(43 downto 30);
row31 <= buf(44 downto 31);
row32 <= buf(45 downto 32);
row33 <= buf(46 downto 33);
row34 <= buf(47 downto 34);
row35 <= buf(48 downto 35);
row36 <= buf(49 downto 36);
row37 <= buf(50 downto 37);
row38 <= buf(51 downto 38);
row39 <= buf(52 downto 39);
row40 <= buf(53 downto 40);
row41 <= buf(54 downto 41);
row42 <= buf(55 downto 42);
row43 <= buf(56 downto 43);
row44 <= buf(57 downto 44);
row45 <= buf(58 downto 45);
row46 <= buf(59 downto 46);
row47 <= buf(60 downto 47);
row48 <= buf(61 downto 48);
row49 <= buf(62 downto 49);
row50 <= buf(63 downto 50);
row51 <= buf(64 downto 51);
row52 <= buf(65 downto 52);
row53 <= buf(66 downto 53);
row54 <= buf(67 downto 54);
row55 <= buf(68 downto 55);
row56 <= buf(69 downto 56);
row57 <= buf(70 downto 57);
row58 <= buf(71 downto 58);
row59 <= buf(72 downto 59);
row60 <= buf(73 downto 60);
row61 <= buf(74 downto 61);
row62 <= buf(75 downto 62);
row63 <= buf(76 downto 63);
row64 <= buf(77 downto 64);
row65 <= buf(78 downto 65);
row66 <= buf(79 downto 66);
row67 <= buf(80 downto 67);
row68 <= buf(81 downto 68);
row69 <= buf(82 downto 69);
row70 <= buf(83 downto 70);
row71 <= buf(84 downto 71);
row72 <= buf(85 downto 72);
row73 <= buf(86 downto 73);
row74 <= buf(87 downto 74);
row75 <= buf(88 downto 75);
row76 <= buf(89 downto 76);
row77 <= buf(90 downto 77);
row78 <= buf(91 downto 78);
row79 <= buf(92 downto 79);
row80 <= buf(93 downto 80);
row81 <= buf(94 downto 81);
row82 <= buf(95 downto 82);
row83 <= buf(96 downto 83);
row84 <= buf(97 downto 84);
row85 <= buf(98 downto 85);
row86 <= buf(99 downto 86);
row87 <= buf(100 downto 87);
row88 <= buf(101 downto 88);
row89 <= buf(102 downto 89);
row90 <= buf(103 downto 90);
row91 <= buf(104 downto 91);
row92 <= buf(105 downto 92);
row93 <= buf(106 downto 93);
row94 <= buf(107 downto 94);
row95 <= buf(108 downto 95);
row96 <= buf(109 downto 96);
row97 <= buf(110 downto 97);
row98 <= buf(111 downto 98);
    end if;
end process dummy_proc;

end architecture behavioral;
